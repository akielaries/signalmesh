/*
 * PLL Example for Gowin FPGAs
 *
 * This module demonstrates how to instantiate a Phase-Locked Loop (PLL)
 * to multiply a clock frequency.
 *
 * IMPORTANT: This is a generic example. For a real design, you should use
 * the Gowin IP Core Generator tool in the Gowin EDA to generate a PLL
 * with parameters validated for your specific device and frequency plan.
 * The tool will provide a customized instantiation template.
 *
 */

module pll_example (
  // --- Inputs ---
  input bank1_3v3_xtal_in, // Input clock from the crystal oscillator (27 MHz)
  input bank3_1v8_sys_rst,      // Active-low reset

  // --- Outputs ---
  output clk_108mhz_out, // Synthesized, faster clock (108 MHz)
  output pll_locked      // High when the PLL output clock is stable
);

wire clk;
wire rst_n;
wire clk_108mhz_internal; // Internal wire for PLL output and feedback

assign clk = bank1_3v3_xtal_in;

assign rst_n = bank3_1v8_sys_rst;
assign clk_108mhz_out = clk_108mhz_internal; // Assign internal wire to output port


// --- PLL Instantiation ---
// The module name (e.g., Gowin_rPLL) and parameters should ideally be
// generated by the Gowin IP Core Generator.
//
// Frequency Calculation:
// F_out = F_in * (FBDIV_SEL / IDIV_SEL) / ODIV_SEL
// 108 MHz = 27 MHz * (20 / 1) / 5
//
// The internal VCO frequency will be:
// F_vco = F_in * (FBDIV_SEL / IDIV_SEL) = 27 * (20 / 1) = 540 MHz
// This VCO frequency is then divided by ODIV_SEL to get the final output.
// A VCO frequency between 400-1600 MHz is typical.

rPLL #(
  .FCLKIN("27"),      // Input clock frequency in MHz
  .IDIV_SEL(0),       // Input Divider (VCO pre-divider)
  .FBDIV_SEL(3),     // Feedback Divider (VCO multiplier)
  .ODIV_SEL(4)        // Output Divider
)
rpll_inst (
  // --- Port Connections ---
  .CLKIN(clk),   // Connect to the 27 MHz input clock
  .RESET(rst_n),         // Connect to the system reset

  .CLKOUT(clk_108mhz_internal), // The generated 108 MHz clock
  .LOCK(pll_locked),      // The PLL lock signal

  // Unused ports can be left blank
  .CLKOUTP(),
  .CLKOUTD(),
  .CLKFB(clk_108mhz_internal), // Explicitly close the feedback loop
  .PSDA(),
  .DUTYDA()
);

endmodule
